// `include "sbox/blind.vh"
// localparam blind_n_rnd = _blind_nrnd(d);
// localparam bcoeff = _bcoeff(d);

// localparam n_random_z = d*(d-1);
// localparam rnd_busz = coeff*n_random_z;
// localparam rnd_busb = bcoeff*blind_n_rnd;

localparam rnd_busz = 2;
localparam rnd_busb = 2;
